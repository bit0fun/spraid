module dump();
	initial begin
		$dumpfile("pload_shift.vcd");
		$dumpvars(0, pload_shift);
		#1;
	end
endmodule
